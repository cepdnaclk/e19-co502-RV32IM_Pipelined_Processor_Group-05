../design/rv32i_decoder_header.vh